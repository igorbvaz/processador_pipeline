module teste(in, out);

input in;
output out;

endmodule