module instruction_memory(endereco, instrucao);

input [31:0] endereco;
output reg [31:0] instrucao;
reg [31:0] instrucoes[31:0];

always @(endereco)
begin
 instrucao=instrucoes[endereco];
end

initial
begin
	instrucoes[0] 	= 32'b11111111111111111111111111111111; //LW
	instrucoes[1] 	= 32'b00111000000100000000000000000011; //SW
	instrucoes[2] 	= 32'b11111111111111111111111111111111; //ADD
	instrucoes[3] 	= 32'b11111111111111111111111111111111; //SUB
	instrucoes[4] 	= 32'b11111111111111111111111111111111; //MUL
	instrucoes[5] 	= 32'b11111111111111111111111111111111; //DIV
	instrucoes[6] 	= 32'b11111111111111111111111111111111; //AND
	instrucoes[7] 	= 32'b11111111111111111111111111111111; //OR
	instrucoes[8] 	= 32'b11111111111111111111111111111111; //SHL
	instrucoes[9] 	= 32'b11111111111111111111111111111111; //SHR
	instrucoes[10] = 32'b11111111111111111111111111111111; //CMP
	instrucoes[11] = 32'b11111111111111111111111111111111; //NOT
	instrucoes[12] = 32'b11111111111111111111111111111111; //JR
	instrucoes[13] = 32'b11111111111111111111111111111111; //JPC
	instrucoes[14] = 32'b11111111111111111111111111111111; //BRFL
	instrucoes[15] = 32'b11111111111111111111111111111111; //CALL
	instrucoes[16] = 32'b11111111111111111111111111111111; //RET
	instrucoes[17] = 32'b11111111111111111111111111111111; //NOP
end

endmodule