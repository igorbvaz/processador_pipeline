module banco_registradores();
endmodule